LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

entity tFlipFlop is
	port(
	
		i_t : in std_logic;
		i_clock : in std_logic;
		o_q, o_qBar : out std_logic

	);
end entity tFlipFlop;

architecture rtl of tFlipFlop is

    begin 


end rtl; 